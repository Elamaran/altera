
module top (
input wire clk, 
input wire rstn,
output wire led[2:0]);

